* D:\Analog_VLSI\eSIM\FOSSEE\eSim\library\SubcircuitLibrary\6T_RAM_sub_ckt\6T_RAM_sub_ckt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/02/22 22:28:02

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M3-Pad1_ Net-_M1-Pad1_ Net-_M2-Pad1_ Net-_M3-Pad1_ mosfet_p		
M5  Net-_M3-Pad1_ Net-_M2-Pad1_ Net-_M1-Pad1_ Net-_M3-Pad1_ mosfet_p		
M2  Net-_M2-Pad1_ Net-_M1-Pad1_ GND GND mosfet_n		
M4  Net-_M1-Pad1_ Net-_M2-Pad1_ GND GND mosfet_n		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ GND mosfet_n		
M6  Net-_M6-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad1_ GND mosfet_n		
U1  Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M6-Pad1_ Net-_M1-Pad1_ PORT		
v1  Net-_M3-Pad1_ GND DC		

.end
