* D:\Analog_VLSI\eSIM\FOSSEE\eSim\library\SubcircuitLibrary\1-bit_RAM_sub_ckt\1-bit_RAM_sub_ckt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/03/22 11:16:26

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
x1  Net-_U2-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ Net-_M1-Pad2_ 6T_RAM_cell		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ writer_ckt		
U4  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U4-Pad3_ Net-_U4-Pad4_ dac_bridge_2		
U3  Net-_U2-Pad2_ Net-_U2-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M4  Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M2  Net-_M1-Pad3_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_n		
M3  Net-_M2-Pad3_ Net-_M3-Pad2_ GND GND mosfet_n		
v1  Net-_M1-Pad1_ GND DC		
M6  Net-_M1-Pad1_ Net-_M1-Pad3_ Net-_M5-Pad1_ Net-_M1-Pad1_ mosfet_p		
M5  Net-_M5-Pad1_ Net-_M1-Pad3_ GND GND mosfet_n		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_M3-Pad2_ Net-_M5-Pad1_ PORT		

.end
